/*------------------------------------------------------------------------------
 * File          : clk_gen.sv
 * Project       : MLProject
 * Author        : epedlh
 * Creation date : Aug 21, 2019
 * Description   :
 *------------------------------------------------------------------------------*/

module clk_gen #() ();


	
endmodule : clk_gen