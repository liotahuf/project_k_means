/*------------------------------------------------------------------------------
 * File          : classify_block_pipe3.sv
 * Project       : MLProject
 * Author        : epedlh
 * Creation date : Oct 27, 2019
 * Description   :
 *------------------------------------------------------------------------------*/

module classify_block_pipe3 #() ();

endmodule : classify_block_pipe3