/*------------------------------------------------------------------------------
 * File          : yyyyyy.sv
 * Project       : MLProject
 * Author        : epedlh
 * Creation date : Jan 12, 2020
 * Description   :
 *------------------------------------------------------------------------------*/

module yyyyyy #() ();



endmodule : yyyyyy