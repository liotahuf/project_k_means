/*------------------------------------------------------------------------------
 * File          : tb_controller.sv
 * Project       : MLProject
 * Author        : epedlh
 * Creation date : Jan 5, 2020
 * Description   :
 *------------------------------------------------------------------------------*/

module tb_controller #() ();

endmodule : tb_controller